-- Copyright (C) 2018  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details.

-- PROGRAM		"Quartus Prime"
-- VERSION		"Version 18.0.0 Build 614 04/24/2018 SJ Lite Edition"
-- CREATED		"Tue May 14 20:33:46 2019"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY fpga IS 
	PORT
	(
		SYSRST :  IN  STD_LOGIC;
		CLK :  IN  STD_LOGIC;
		SLIDERS :  IN  STD_LOGIC_VECTOR(9 DOWNTO 0);
		PCSRC :  OUT  STD_LOGIC;
		PCWR :  OUT  STD_LOGIC;
		REGDST :  OUT  STD_LOGIC;
		REGWR :  OUT  STD_LOGIC;
		ALUSRCB :  OUT  STD_LOGIC;
		CPSRWR :  OUT  STD_LOGIC;
		MEMRD :  OUT  STD_LOGIC;
		MEMWR :  OUT  STD_LOGIC;
		MULTIPLY :  OUT  STD_LOGIC;
		RDORBL :  OUT  STD_LOGIC;
		PCLRBR :  OUT  STD_LOGIC;
		C :  OUT  STD_LOGIC;
		V :  OUT  STD_LOGIC;
		N :  OUT  STD_LOGIC;
		Z :  OUT  STD_LOGIC;
		ALUS :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		BRADDR :  OUT  STD_LOGIC_VECTOR(31 DOWNTO 0);
		EXTS :  OUT  STD_LOGIC_VECTOR(1 DOWNTO 0);
		INSTR :  OUT  STD_LOGIC_VECTOR(31 DOWNTO 0);
		LEDS :  OUT  STD_LOGIC_VECTOR(9 DOWNTO 0);
		PC4 :  OUT  STD_LOGIC_VECTOR(31 DOWNTO 0);
		REGSRC :  OUT  STD_LOGIC_VECTOR(1 DOWNTO 0);
		ROTATE :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		SEG0 :  OUT  STD_LOGIC_VECTOR(7 DOWNTO 0);
		SEG1 :  OUT  STD_LOGIC_VECTOR(7 DOWNTO 0);
		SEG2 :  OUT  STD_LOGIC_VECTOR(7 DOWNTO 0);
		SEG3 :  OUT  STD_LOGIC_VECTOR(7 DOWNTO 0);
		SEG4 :  OUT  STD_LOGIC_VECTOR(7 DOWNTO 0);
		SEG5 :  OUT  STD_LOGIC_VECTOR(7 DOWNTO 0);
		WB :  OUT  STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END fpga;

ARCHITECTURE bdf_type OF fpga IS 

COMPONENT spc
	PORT(RST : IN STD_LOGIC;
		 CLK : IN STD_LOGIC;
		 MEMDATAIN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 PCSRC : OUT STD_LOGIC;
		 PCWR : OUT STD_LOGIC;
		 REGDST : OUT STD_LOGIC;
		 REGWR : OUT STD_LOGIC;
		 ALUSRCB : OUT STD_LOGIC;
		 CPSRWR : OUT STD_LOGIC;
		 MEMRD : OUT STD_LOGIC;
		 MEMWR : OUT STD_LOGIC;
		 MULTIPLY : OUT STD_LOGIC;
		 RDORBL : OUT STD_LOGIC;
		 PCLRBR : OUT STD_LOGIC;
		 C : OUT STD_LOGIC;
		 V : OUT STD_LOGIC;
		 N : OUT STD_LOGIC;
		 Z : OUT STD_LOGIC;
		 ALUS : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 BRADDR : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 EXTS : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		 INSTR : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 MEMADDR : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 MEMDATAOUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 PC4 : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 REGSRC : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		 ROTATE : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 WB : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT dmem
	PORT(MEMWR : IN STD_LOGIC;
		 RST : IN STD_LOGIC;
		 CLK : IN STD_LOGIC;
		 A : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 WD : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 RD : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT busmux2to1
	PORT(S : IN STD_LOGIC;
		 D0 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 D1 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Y : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT synchronizer
	PORT(SYSRST : IN STD_LOGIC;
		 CLK : IN STD_LOGIC;
		 RST : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT reg10
	PORT(LD : IN STD_LOGIC;
		 RST : IN STD_LOGIC;
		 CLK : IN STD_LOGIC;
		 D : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
		 Q : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT led
	PORT(LD : IN STD_LOGIC;
		 RST : IN STD_LOGIC;
		 CLK : IN STD_LOGIC;
		 D : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Q : OUT STD_LOGIC_VECTOR(9 DOWNTO 0)
	);
END COMPONENT;

COMPONENT seg7decode
	PORT(LD : IN STD_LOGIC;
		 RST : IN STD_LOGIC;
		 CLK : IN STD_LOGIC;
		 INP : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 SEG0 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 SEG1 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 SEG2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 SEG3 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 SEG4 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 SEG5 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT addressdecoder
	PORT(MEMRD : IN STD_LOGIC;
		 MEMWR : IN STD_LOGIC;
		 ADDR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 LD2 : OUT STD_LOGIC;
		 LD1 : OUT STD_LOGIC;
		 LD0 : OUT STD_LOGIC;
		 DATAS : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL	DATAS :  STD_LOGIC;
SIGNAL	LD0 :  STD_LOGIC;
SIGNAL	LD1 :  STD_LOGIC;
SIGNAL	LD2 :  STD_LOGIC;
SIGNAL	MEMRD_ALTERA_SYNTHESIZED :  STD_LOGIC;
SIGNAL	MEMWR_ALTERA_SYNTHESIZED :  STD_LOGIC;
SIGNAL	RST :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;


BEGIN 
SYNTHESIZED_WIRE_5 <= '1';



b2v_inst : spc
PORT MAP(RST => RST,
		 CLK => CLK,
		 MEMDATAIN => SYNTHESIZED_WIRE_0,
		 PCSRC => PCSRC,
		 PCWR => PCWR,
		 REGDST => REGDST,
		 REGWR => REGWR,
		 ALUSRCB => ALUSRCB,
		 CPSRWR => CPSRWR,
		 MEMRD => MEMRD_ALTERA_SYNTHESIZED,
		 MEMWR => MEMWR_ALTERA_SYNTHESIZED,
		 MULTIPLY => MULTIPLY,
		 RDORBL => RDORBL,
		 PCLRBR => PCLRBR,
		 C => C,
		 V => V,
		 N => N,
		 Z => Z,
		 ALUS => ALUS,
		 BRADDR => BRADDR,
		 EXTS => EXTS,
		 INSTR => INSTR,
		 MEMADDR => SYNTHESIZED_WIRE_9,
		 MEMDATAOUT => SYNTHESIZED_WIRE_10,
		 PC4 => PC4,
		 REGSRC => REGSRC,
		 ROTATE => ROTATE,
		 WB => WB);


b2v_inst1 : dmem
PORT MAP(MEMWR => LD2,
		 RST => RST,
		 CLK => CLK,
		 A => SYNTHESIZED_WIRE_9,
		 WD => SYNTHESIZED_WIRE_10,
		 RD => SYNTHESIZED_WIRE_4);


b2v_inst2 : busmux2to1
PORT MAP(S => DATAS,
		 D0 => SYNTHESIZED_WIRE_3,
		 D1 => SYNTHESIZED_WIRE_4,
		 Y => SYNTHESIZED_WIRE_0);


b2v_inst3 : synchronizer
PORT MAP(SYSRST => SYSRST,
		 CLK => CLK,
		 RST => RST);


b2v_inst4 : reg10
PORT MAP(LD => SYNTHESIZED_WIRE_5,
		 RST => RST,
		 CLK => CLK,
		 D => SLIDERS,
		 Q => SYNTHESIZED_WIRE_3);



b2v_inst7 : led
PORT MAP(LD => LD1,
		 RST => RST,
		 CLK => CLK,
		 D => SYNTHESIZED_WIRE_10,
		 Q => LEDS);


b2v_inst8 : seg7decode
PORT MAP(LD => LD0,
		 RST => RST,
		 CLK => CLK,
		 INP => SYNTHESIZED_WIRE_10,
		 SEG0 => SEG0,
		 SEG1 => SEG1,
		 SEG2 => SEG2,
		 SEG3 => SEG3,
		 SEG4 => SEG4,
		 SEG5 => SEG5);


b2v_inst9 : addressdecoder
PORT MAP(MEMRD => MEMRD_ALTERA_SYNTHESIZED,
		 MEMWR => MEMWR_ALTERA_SYNTHESIZED,
		 ADDR => SYNTHESIZED_WIRE_9,
		 LD2 => LD2,
		 LD1 => LD1,
		 LD0 => LD0,
		 DATAS => DATAS);

MEMRD <= MEMRD_ALTERA_SYNTHESIZED;
MEMWR <= MEMWR_ALTERA_SYNTHESIZED;

END bdf_type;